
module unsaved (
	clk_clk,
	pll_clk_50mhz_clk,
	reset_reset_n);	

	input		clk_clk;
	output		pll_clk_50mhz_clk;
	input		reset_reset_n;
endmodule
