
module InternalClock (
	oscena,
	clkout);	

	input		oscena;
	output		clkout;
endmodule
